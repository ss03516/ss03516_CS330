library verilog;
use verilog.vl_types.all;
entity MUX is
    port(
        a               : in     vl_logic_vector(63 downto 0);
        b               : in     vl_logic_vector(63 downto 0);
        \select\        : in     vl_logic;
        data            : out    vl_logic_vector(63 downto 0)
    );
end MUX;
